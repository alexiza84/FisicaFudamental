��  CCircuit��  CSerializeHack           ��  CPart              ���  CECapacitor��  CValue  3Q[_    100�F(    ,C��6?      �?�F �� 	 CTerminal  h8iM         L            �  �  hdiy                            \Ltd        ��             �� 
 CVoltmeter��  CMeter  �Y�g     0.00(    �  �@�U         L                �  �l��                             �T�l        ��      ��  CSPDT��  CToggle   8 X         �  (1)        L               �  � !            "@          �  �01        L            �    4          ��    �� 	 CResistor
�  �q�    6k          p�@      �?k  �  �X�m         L               �  ����                       �    �l��         ��      �
�  p�$    58k        R�@      �?k  �  �(�)            "@          �  `(u)            "@            t$�,    #    ��      ��  CBattery
�  +qS    9V(         "@      �? V �  `Xam             "@          �  `�a�                            Tll�     (    ��                    ���  CWire  h8�9      +�  �8�A       +�  0(i)      +�  `(aY       +�  h�i�        +�  hxi�        +�  h���       +�  h(i9       +�  � �)       +�  �(�)      +�  �0�Y       +�  �0�1      +�  `���       +�  ��i�                     �                             3    1  -    2   .  4   7   6      9 # # 5 $ / $ ( / ( ) ) 8  - ,   3 $ ( 1 9  2 0  . ,  5 # 4 7  6  )   8 0   &        �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 