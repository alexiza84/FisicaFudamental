��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � B�     
Resistor 5      �  Q�'    
Resistor 6      �  �9
G    
Resistor 8      �  1B?    
Resistor 4      �  	H    Resistor 10      �  �� ��     
Resistor 9      �  iBw    
Resistor 3      �  �� �     
Resistor 2      �  �� ��     
Resistor 1      �  �i�w    
Resistor 7                    ���  CLED_G�� 	 CTerminal  Pe         �0z��@���&|i?  �  |�        �|j:�@���&|i�    d$|        ��      ��  �P�e         �0z��@ ��&|i?  �  �|��        �|j:�@ ��&|i�    �d�|        ��      ��  L a!        �2�ď @ ��&|i?  �    5!                  ��&|i�    4L4       ��      ��  L a        �2�ď @ ��&|i?  �    5                  ��&|i�    4�L       ��      ��  L�a�        �2�ď @ ��&|i?  �   �5�                  ��&|i�    4�L�    "   ��      ��  L�a�        �2�ď @ ��&|i?  �   �5�                  ��&|i�    4�L�    %   ��      ��  CSPST��  CToggle  �(�      (   �   ��        �2�ď @          �   ��         �0z��@            ���    +      ��    '�)�  X x@     -   �  P<QQ     	        "@h��&|�?  �  PQ%              "@h��&|��    L$T<    /     ��    �� 	 CResistor��  CValue  �$    1         �?      �?   �  (!)        �0z��@ ��&|��  �  �(�)        �{���@ ��&|�?    �$,    5    ��      1�3�  X.x<    1         �?      �?   �  t@�A        ��>���@ ��&|��  �  H@]A        _�����@ ��&|�?    \<tD    9    ��      1�3�  �F�T    1         �?      �?   �  �X�Y        �{���@ ��o�p�  �  �X�Y        ��>���@ ��o�p?    �T�\    =    ��      1�3�  ��,    1         �?      �?   �  �0�1        �{���@ ��o�p�  �  �0�1        ��>���@ ��o�p?    �,�4    A    ��      1�3�  �� �    1         �?      �?   �  ��	        �{���@ ��o�p�  �  ��	        ��>���@ ��o�p?    ��    E    ��      1�3�  �� �    220        �k@      �?   �  ��        7�k�@h��&|��  �  ��             "@h��&|�?    ��    I    ��      1�3�  �� �    1         �?      �?   �  �	     
   NEMX��@ ��&|��  �  ��      	 7�k�@ ��&|�?    ��    M    ��      ��  CBattery3�  iCw    9V(          "@      �? V �  PPQe      	 	       "@h��&|��  �  P|Q�                h��&|�?    Dd\|     R    ��      1�3�  F8T    1         �?      �?   �  4XIY        _�����@ ��o�p�  �  XY     
   NEMX��@ ��o�p?    T4\    V    ��      1�3�  � 8    1         �?      �?   �  4I	        _�����@ ��o�p�  �  	     
   NEMX��@ ��o�p?    4    Z    ��      1�3�  8$    1         �?      �?   �  4(I)        _�����@ ��o�p�  �  ()     
   NEMX��@ ��o�p?    $4,    ^    ��      ��  �P�e         �0z��@���&|i?  �  �|��        �|j:�@���&|i�    �d�|     a   ��      ��  �P�e         �0z��@���&|i?  �  �|��        �|j:�@���&|i�    �d�|     d   ��      '�)�  x���      f   �  p�q�        �|j:�@          �  ppq�         �0z��@            l�t�    h      ��    ��  T�i�        �|j:�@@��o�p?  �  (�=�        �2�ď @@��o�p�    <�T�    k   ��      ��  T�i�        �|j:�@���o�p?  �  (�=�        �2�ď @���o�p�    <�T�    n   ��      ��  T�i�        �|j:�@ ��o�p?  �  (�=�        �2�ď @ ��o�p�    <�T    q   ��                    ���  CWire  `�a�       t�  `�a�       t�  `��      t�  �PQ      t�  ���      t�  �P�Q      t�  ����      t�   �!        t�   �!�        t�  P�!�       t�  P�Q�        t�  h�i�       t�    !!        t�  ` a!       t�  `�a       t�   �!�        t�  (�)�       t�  (�)�       t�   �)�      t�  0 q!      t�    1!      t�  0 1a       t�   `1a      t�   `�       t�  P�      t�  (�)�       t�  p�q�       t�  p���      t�  ����       t�  ����      t�  ����      t�    !)       t�  �(�1       t�  ��)       t�  �(�)      t�  �0�Y       t�  p qq       t�  �@�Y       t�  �0�A       t�  �@�A      t�  ��1       t�  H(IA       t�  H@IY       t�  	      
 t�  	)      
 t�  (	Y      
 t�  HI)       t�  �P�Q      t�  �P�Q      t�  � �Q       t�  p �!      t�  h�i�       t�  h�i�       t�  h�q�                    �                             x    y  z    {   �  �    �   |   " " v # � # % % u & � & + + � , � , / / R 0 � 0 5 5 � 6 � 6 9 9 � : � : = = � > � > A A � B � B E E � F � F I I N J � J M M � N I N R / R S S  V V � W � W Z Z � [ � [ ^ ^ � _ � _ a � a b b � d � d e e � h h � i � i k k � l � l n n � o � o q q � r � r v � " w u +     a x b y } � & ~  | S ~ k q      % � # } � � o � w � � � � � � � � � � , 0 J l r h � � � � � e � � { � 5 � � E � � 6 A = � i � > B � 9 � F � ^ : � V [ M � � _ W Z � � z d � � � � � n � � � � �   P         �4s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 