��  CCircuit��  CSerializeHack           ��  CPart              ���  CECapacitor��  CValue  3Q[_    100�F(    -C��6?      �?�F �� 	 CTerminal  h8iM         P�*w�ƕ>P��_����  �  hdiy                 P��_���=    \Ltd        ��      M��_���=��  CSPDT��  CToggle   8 X         �  (1)        P�*w�ƕ>M��_���=  �  � !            "@          �  �01        P�*w�ƕ>M��_����    4          ��    �� 	 CResistor
�  �q�    10k          ��@      �?k  �  �X�m         P�*w�ƕ>M��_���=  �  ����                 M��_����    �l��         ��      �
�  p�$    10k        ��@      �?k  �  �(�)            "@          �  `(u)            "@            t$�,        ��      �� 
 CVoltmeter��  CMeter  �Q�_     0.32(    �  �8�M         P�*w�ƕ>          �  �d�y                             �L�d     #   ��      ��  CBattery
�  +qS    9V(         "@      �? V �  `Xam             "@          �  `�a�                            Tll�     (    ��                    ���  CWire  � �)       +�  �(�)      +�  �0�Y       +�  �0�1      +�  0(i)      +�  `���       +�  ��i�       +�  `(aY       +�  h(i9       +�  h(�)      +�  �(�9       +�  h���       +�  �x��        +�  hxi�                      �                             4    9   0  ,   /   .    2   -  3  # 6 # $ $ 8 ( 3 ( ) ) 1  -  , /  .   4 )  1 9  ( 5  0 6 5 # 2 8 $ 7  7   &        �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 