��  CCircuit��  CSerializeHack           ��  CPart              ���  CNPN��  CDummyValue  p�p�    100hFE            Y@      �? hFE �� 	 CTerminal  p�q�         �M=�ͼ@Fs4볪}?  �  H�]�        ���o���?��h��?  �  p�q�                 ��Ԉ��}�    \�x�         ��      �� 	 CResistor��  CValue  �(�    1k        @�@      �?k  �  $�9�        ���o���?ɖh���  �  � ��        �B5����?ɖh��?    �$�        ��      ��  � 	�     10k          ��@      �?k  �  � ��          �B5����?J�:S�?  �  � � 1                 J�:S��    � �          ��      ��  � �� �    10k          ��@      �?k  �  � p� �         �M=�ͼ@详9�F#?  �  � �� �        �B5����?详9�F#�    � �� �         ��      ��  CLED�   HI        �M=�ͼ@(J��uUֺ  �  ,HAI        �M=�ͼ@(J��uU�:    <,\         ��      ��  P6pD    600        ��@      �?   �  lH�I        �M=�ͼ@0��b�/f�  �  @HUI      	 �M=�ͼ@0��b�/f<    TDlL    $    ��      �
�  P�P�    100hFE            Y@      �? hFE �  P�Q�         js��4�?������C?  �  (�=�        �JV��?�� �&1?  �  P�Q                 �͙���F�    <�X�     (    ��      ��  ���    1k        @�@      �?k  �  ��        �JV��?�� �&1�  �  ����        �	[��?�� �&1?    ���    -    ��      ��  ��    10k          ��@      �?k  �  ���         �	[��?�ҳGw?  �  �$�9                 �ҳGw�    ��$     1    ��      ��  ����    10k          ��@      �?k  �  �x��         �M=�ͼ@#+j�#?  �  ����        �	[��?#+j�#�    ����     5    ��      ��  �P�Q        �M=�ͼ@ �����C?  �  P!Q        eAk���? �����C�    �Dd    8    ��      ��  0>PL    600        ��@      �?   �  LPaQ        js��4�?������C�  �   P5Q      	 eAk���?������C?    4LLT    <    ��      ��  CBattery�  3 � [ �     9V(          "@      �? V �  h h i }               "@��C�8'��  �  h � i �                 ��C�8'�?    \ | t �      A    ��      ��  p �     600        ��@      �?   �  �  �!         �M=�ͼ@2��{,���  �  `  u!       	 ��G��l@2��{,��?    t �$     E    ��      ��  � p � �          �]�'l�?�����?  �  � � � �                  ������    � � � �      H  
 ��      ��  � p � �          �]�'l�?�����?  �  � � � �                  ������    � � � �      K  
 ��      ��  � p � �          �]�'l�?�����?  �  � � � �                  ������    � � � �      N  
 ��      ��  � 9 � G     220          �k@      �?   �  �   � 5               "@H8*�6��?  �  � L � a         �]�'l�?H8*�6���    � 4 � L      R    ��      ��     5!              "@���{,��?  �  L  a!         ��G��l@���{,���    4 L4     U   ��      ��  � a o     10k          ��@      �?k  �  H ]               "@��H�}M?  �  t �                  ��H�}M�    \ t      Y    ��      ��  � � �     10k          ��@      �?k  �  � �                             �  � 	                             � �      ]    ��      ��  (� H�     1k        @�@      �?k  �  D� Y�      
   ?�f_��W>��5M�`�=  �  � -�                  ��5M�`��    ,� D�     a    ��      �
�  �� ��     100hFE            Y@      �? hFE �  �� ��          �M=�ͼ@�-�ϬH�=  �  h� }�      
   ?�f_��W>��5M�`��  �  �� ��                  �%y޽    |� ��      e    ��      �
�  �� ��     100hFE            Y@      �? hFE �  �� ��          ��{��,@!G Ƿ>  �  �� ��         �Z9�2�?��Ѳ�y=  �  �� ��                  �^�l@��    �� ��      j    ��      ��  @� `�     1k        @�@      �?k  �  \� q�         �Z9�2�?��T����  �  0� E�      	   w�4�3�?��T����=    D� \�     o    ��      ��  � +�     10k          ��@      �?k  �  0� 1�       	   w�4�3�?rXG���>  �  0� 1                 rXG����    ,� 4�      s    ��      ��   �  �     1.6M        j8A      �?M  �  � 1�      	   w�4�3�?k$a���  �  �� �         �M=�ͼ@k$a��>    � �     w    ��      ��  �6  D     600        ��@      �?   �  �H I                  ��<��  �  �H �I       	 z��È?�>��<��=    �D �L     {    ��      ��  �H �I         �Z9�2�?��<��=  �  �H �I         z��È?�>��<��    �< �\     ~    ��      ��  8  M!       	 ��/3ͼ@�G Ƿ>  �  d  y!         ��{��,@�G Ƿ�    L d4     �    ��      ��   (     600        ��@      �?   �  $  9!         ��/3ͼ@�6 Ƿ�  �  �  !         �M=�ͼ@�6 Ƿ>     $$     �    ��                    ���  CWire  � H� q       ��  �  � I       ��  �  �!      ���� 
 CCrossOver  ��        �  �!       ��  � �I       ��  ��       ��  0�       ��  ��9        ��  P8�9       ��  p�q1        ��  p0q9        ��  p8�9       ��  �8Q9       ��  �P�Q      ��  �H�Q       ��  �H�I      ��  �H�I      ��  �  �!       ����  ��        �1       ��  �  �!       ��  � 0q1       ��  p���      ��  8�I�      ��  � �� �       ��  � �� �       ��  � HI      ��  P�a�      ��  `Pa�       ��  P Q9        ��  �)�      ��  ����       ��  ����       ��  �P�y       ��  �H��       ��  � p � q       ��  � ` � a       ��  � ` � q        ��  � p � q       ��  � p � q       ��  � � � �        ��  � � � �        ��  � � � �        ��  � � � �         ��  h � i �         ��  h   � !       ��  h   i i        ��    I        ��    !!       ��  h � � �        ��  � � �        ��  � � � �        ��  � � � 	        ��  � 	       ��  � �         ��  � �         ��  X� i�      
 ��  �� �	        ��  �  ��        ��  �� ��       ��  ��        ��  �	       ��  0� 1�       	 ��  0� 1�       	 ��  �  ��        ��  xH �I       ��  p� y�       ��  x� ��       ��  H         ��  �       ��  �� �        ��  �� ��       ��  �� ��        ����  v� |�         xH y�        ����  v� |�         8� ��       ��  x  yA        ��  8@ yA       ��  8@ 9�        ��  �  �!       ��  �   !                     �                             �   �    �   �  �   �    �  �    �   �   ! ! % $ $ � % ! % ( � ( ) � ) * * � - - � . � . 1 � 1 2 2 � 5 � 5 6 6 � 8 � 8 9 9 = < < � = 9 = A � A B B � E E � F V F H � H I I � K � K L L � N � N O O � R � R S S � U � U V V F Y � Y Z Z � ] � ] ^ ^ � a a � b � b e � e f � f g g � j � j k � k l l � o o � p � p s � s t t � w w � x � x { { � |  | ~ � ~   | � � � � � � � � � � � � �  � � � � � � � � � � � � � � � � � �  � � � � 2 � � � 8 � � � � $ � � � � � � t � �  �  �     �  �   ( � < � * � - ) 6 . � 1 � 5 � � H K � S � � N � � � O I � L � � � � B � � R � A � Y � U � � � � � � � � � � � ] Z b a f g � E � e � � � ^ � � s w p � x � ~ o � � k { � � � l � � j � � � � � � � � � � � � � � � � � � � �   ?         �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 